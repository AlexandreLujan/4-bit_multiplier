PACKAGE MyPackage IS

	COMPONENT ADDER
	PORT (
		A, B, C_IN : IN BIT;
		C_OUT, S   : OUT BIT
	);
	END COMPONENT;
	
	COMPONENT TOP_BLOCK
	PORT (        
		MK, MK1, Q0, Q1, CIN : IN BIT;
		COUT, SI   				: OUT BIT
	);
	END COMPONENT;
	
	COMPONENT BOTTOM_BLOCK
	PORT (        
		MK, PPI, QJ, CIN 	: IN BIT;
		COUT, SI   			: OUT BIT
	);
	END COMPONENT;
	
	COMPONENT MULTIPLIER 
   PORT (
		M, Q : IN  BIT_VECTOR (3 DOWNTO 0);
		P     : OUT BIT_VECTOR (7 DOWNTO 0)
	);
	END COMPONENT;
	   
END MyPackage;

PACKAGE BODY MyPackage IS
	CONSTANT CONSTANTE_GLOBAL: INTEGER := 200;
END MyPackage;