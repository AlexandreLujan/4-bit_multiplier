LIBRARY work;
USE work.MyPackage.all;

ENTITY TESTBENCH IS
END ENTITY;

ARCHITECTURE RTL OF TESTBENCH IS

	SIGNAL S_M, S_Q : BIT_VECTOR (3 DOWNTO 0);
	SIGNAL S_P: BIT_VECTOR (7 DOWNTO 0);
	
BEGIN

    MULTIPLIER_0 : MULTIPLIER
		PORT MAP (
			M   => S_M,
			Q   => S_Q,
			P   => S_P
		);
	
	S_M <= "0010" AFTER 0ns, "1111" AFTER 40ns;
	S_Q <= "0110" AFTER 0ns, "1111" AFTER 40ns;
		  
END ARCHITECTURE;